.title KiCad schematic
V1 Net-_R1-Pad1_ GND dc 5
R1 Net-_R1-Pad1_ Net-_C1-Pad1_ 10
C1 Net-_C1-Pad1_ GND 50U
R2 Net-_C1-Pad1_ GND 1M
.TRAN 5u 1 
.end
